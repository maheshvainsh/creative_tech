package pcie_rc_pkg;
import uvm_pkg::*;//compile uvm lib
`include "uvm_macros.svh"
`include "pcie_rc_monitor.sv"
`include "pcie_rc_driver.sv"
`include "pcie_rc_sequencer.sv"
`include "pcie_rc_agent.sv"
endpackage : pcie_rc_pkg
