package pcie_sw_pkg;
import uvm_pkg::*;//compile uvm lib
`include "uvm_macros.svh"
`include "pcie_sw_monitor.sv"
`include "pcie_sw_driver.sv"
`include "pcie_sw_sequencer.sv"

`include "pcie_sw_agent.sv"
endpackage : pcie_sw_pkg
