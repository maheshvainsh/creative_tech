//----------------------------------------------------------------------
// Project       : AUURORALANE
// File          : pcie_test_lib.sv
//----------------------------------------------------------------------
// Created by    : MAHESH VANISH
//               : RUTVIK MAKWANA
// Creation Date : 2025-09-06
//----------------------------------------------------------------------
// Description   : 
//                 
//----------------------------------------------------------------------
`ifndef PCIE_TEST_LIB_SV
`define PCIE_TEST_LIB_SV

`include "pcie_base_test.sv"

`endif //PCIE_TEST_LIB_SV
