`ifndef PCIE_PARAMETER_SV
`define PCIE_PARAMETER_SV

//keep define common paramter here
parameter LAN_WIDTH   =1;
parameter DATA_WIDTH = 32;
parameter ADDR_WIDTH = 32;
parameter NO_OF_VC = 3;

`endif //PCIE_PARAMETER_SV
