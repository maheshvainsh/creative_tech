//----------------------------------------------------------------------
// Project       : AUURORALANE
// File          : pcie_ral_pkg.sv
//----------------------------------------------------------------------
// Created by    : MAHESH VANISH
//               : RUTVIK MAKWANA
// Creation Date : 2025-09-06
//----------------------------------------------------------------------
// Description   : 
//                 
//----------------------------------------------------------------------
 `include "pcie_config_reg.sv"
 `include "pcie_cfg_regfile.sv"
 `include "pcie_cfg_block.sv"
 `include "pcie_reg_adapter.sv"
