`ifndef PCIE_SEQ_LIB_SVH
`define PCIE_SEQ_LIB_SVH

`include "pcie_base_sequence.sv"

`endif //PCIE_SEQ_LIB_SVH
