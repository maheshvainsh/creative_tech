
//keep define common paramter here
parameter LAN_WIDTH   =1;
parameter DATA_WIDTH = 32;
parameter ADDR_WIDTH = 32;
parameter NO_OF_VC = 3;
