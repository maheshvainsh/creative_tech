//first progame on git repo
module tb ;



initial begin
$display("HELLO WORLD");

end






endmodule : tb
