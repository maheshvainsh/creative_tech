 `include "pcie_config_reg.sv"
 `include "pcie_cfg_regfile.sv"
 `include "pcie_cfg_block.sv"
 `include "pcie_reg_adapter.sv"
