//----------------------------------------------------------------------
// Project       : AUURORALANE
// File          : pcie_if.sv
//----------------------------------------------------------------------
// Created by    : MAHESH VANISH
//               : RUTVIK MAKWANA
// Creation Date : 2025-09-06
//----------------------------------------------------------------------
// Description   : 
//                 
//----------------------------------------------------------------------
`ifndef PCIE_IF_SV
`define PCIE_IF_SV

interface pcie_if ;

//tx link diff pair 
/*logic tx_p[NUMBER_OF_LANE];
logic tx_n[NUMBER_OF_LANE];

//rx link with diff pair
logic tx_p[NUMBER_OF_LANE];
logic tx_n[NUMBER_OF_LANE];*/


endinterface : pcie_if
`endif //PCIE_IF_SV
