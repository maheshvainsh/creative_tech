`ifndef PCIE_TEST_LIB_SV
`define PCIE_TEST_LIB_SV

`include "pcie_base_test.sv"

`endif //PCIE_TEST_LIB_SV
