//----------------------------------------------------------------------
// Project       : AUURORALANE
// File          : pcie_seq_lib.svh
//----------------------------------------------------------------------
// Created by    : MAHESH VANISH
//               : RUTVIK MAKWANA
// Creation Date : 2025-09-06
//----------------------------------------------------------------------
// Description   : 
//                 
//----------------------------------------------------------------------
`ifndef PCIE_SEQ_LIB_SVH
`define PCIE_SEQ_LIB_SVH

`include "pcie_base_sequence.sv"

`endif //PCIE_SEQ_LIB_SVH
