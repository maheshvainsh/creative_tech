package pcie_ep_pkg;
import uvm_pkg::*;//compile uvm lib
`include "uvm_macros.svh"

`include "pcie_ep_monitor.sv"
`include "pcie_ep_driver.sv"
`include "pcie_ep_sequencer.sv"
`include "pcie_ep_agent.sv"

endpackage : pcie_ep_pkg
