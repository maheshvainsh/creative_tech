//classs mem model
//add[]
//data





//write(add, data)

  //writmemh("txt", add,data,byte enable)
//add++





//read(ref data)
//readmemh(data)


//endclass
